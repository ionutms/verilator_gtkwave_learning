module test; // Test module
    initial $display("Hello"); // Display message from the test module
endmodule // End of test module